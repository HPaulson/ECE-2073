    Mac OS X            	   2  G     y    ��������                          ATTR      y  `                   `   �  "com.apple.LaunchServices.OpenWith      �   $  com.apple.decmpfs           com.apple.lastuseddate#PS      *   H  com.apple.macl     r     com.macromates.selectionRange      w     com.macromates.visibleIndex  bplist00�WversionTpath_bundleidentifier _$/Applications/Visual Studio Code.app_com.microsoft.VSCode/1X                            ofpmc  ��         �t�TBT���[:�,aEb    f82     ;2���K��%����                                                      28:8588